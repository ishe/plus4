`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//  Copyright 2013-2016 Istvan Hegedus
//
//  FPGATED is free software: you can redistribute it and/or modify
//  it under the terms of the GNU General Public License as published by
//  the Free Software Foundation, either version 3 of the License, or
//  (at your option) any later version.
//
//  FPGATED is distributed in the hope that it will be useful,
//  but WITHOUT ANY WARRANTY; without even the implied warranty of
//  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//  GNU General Public License for more details.
//
//  You should have received a copy of the GNU General Public License
//  along with this program.  If not, see <http://www.gnu.org/licenses/>. 
//
// 
// Create Date:    12:02:05 16/09/2016 
// Design Name: 	 Commodore Plus 4 in an FPGA
// Module Name:    PLUS4.v
// Project Name: 	 FPGATED Papilio Pro edition
//
// Description: 	
//	This module provides the top level framework for FPGATED. It implements a Commodore Plus 4 computer without expansion port.
// It is written for Papilio FPGATED wing 1.x but can be easily modified for any other platforms.
//
// Revision history: 
// 1.0   16.09.2016			 Commodore Plus 4 shell created, SDRAM based memory (Papilio Pro)
// 1.1	15.12.2016			 Bootstrap function implemented, loads ROMs to SDRAM
//
//	Comments:                This module is based on c16.v which is part of the original FPGATED design and it makes use of Papilio Pro platform's sdram.
//									 Using the sdram of Papilio Pro more ROM can be used thus it is possible to implement a Commodore Plus 4.
//	                         Note however that it is not a complete Plus 4 system; expansion port,user port and ACIA is not yet implemented
//
//////////////////////////////////////////////////////////////////////////////////

module Plus4(
	input wire CLK32,
	input wire RESET,
	output wire HSYNC,
	output wire VSYNC,
	output wire [3:0] RED,
	output wire [3:0] GREEN,
	output wire [3:0] BLUE,
	input PS2DAT,
	input PS2CLK,
	output IEC_DATAOUT,
	input IEC_DATAIN,
	output IEC_CLKOUT,
	input IEC_CLKIN,
	output IEC_ATNOUT,
// input IEC_ATNIN,
	output IEC_RESET,
	output AUDIO_L,
	output AUDIO_R,
//	input RGBS,

	//  SDRAM signals on Papilio Pro board
	output wire [11:0] SDRAM_ADDR,
	inout wire [15:0] SDRAM_DATA,
	output wire SDRAM_DQML,
	output wire SDRAM_DQMH,
	output wire [1:0] SDRAM_BA,
	output wire SDRAM_nWE,
	output wire SDRAM_nCAS,
	output wire SDRAM_nRAS,
	output wire SDRAM_CS,
	output wire SDRAM_CLK,
	output wire SDRAM_CKE,

	// FLASH chip signals on Papilio Pro board
	output wire FLASH_CS,
	output wire FLASH_CK,
	output wire FLASH_SI,
	input wire FLASH_SO
    );

wire CLK28;							// This is the main system clock generated by DCM. It must be 4*dot clk so 28.375152MHz for PAL (1.6*PAL system's clock) and 28.63636 for NTSC (2*NTSC system's clock) 
wire phi0;
reg phi0_prev;
wire [15:0] plus4_addr;
wire [15:0] ted_addr;
wire [15:0] cpu_addr;
wire [15:0] boot_addr;
wire [5:0] boot_addrext;
wire [5:0] plus4_addrext;
wire [7:0] boot_data;
wire [7:0] config_data;
wire [7:0] plus4_data,ted_data,ram_data,cpu_data,port_in,port_out,keyport_data;
wire [7:0] keyboard_row,kbus,key;
wire [7:0] keyscancode;
wire keyreceived;
wire [6:0] plus4_color;
wire mux;
wire cpuenable;
wire aec;
wire rdy;
wire sound;
wire FD0x,FD1x,FD2x,FD3x,FDDx,FD9x;
reg FDDx_prev,FD9x_prev;
wire phi2;
wire KERN;
wire raminitdone;

reg [3:0] romselect=0;						// Plus4/C16 motherboard U21 ROM selector register
reg [3:0] Kernalver=4'h0;					// Kernal ROM alternative version selector 1-16
reg [3:0] Basicver=4'h0;					// Basic ROM alternative version selector 1-16
reg [3:0] FunctionLver=4'h0;				// Function ROM alternative version selector 1-16 (Low)
reg [3:0] FunctionHver=4'h0;				// Function ROM alternative version selector 1-16 (High)
reg [3:0] C1Lver=4'h0;						// Cartridge ROM1 alternative version selector 1-16 (Low)
reg [3:0] C1Hver=4'h0;						// Cartridge ROM1 alternative version selector 1-16 (Low)
reg [3:0] C2Lver=4'h0;						// Cartridge ROM2 alternative version selector 1-16 (Low)
reg [3:0] C2Hver=4'h0;						// Cartridge ROM2 alternative version selector 1-16 (High)
reg [3:0] romversion;						// Addressed ROM's version (1-16)
reg [5:0] romaddrext;						// ROM address extension 4M ROM area (see sdram controller)
reg [5:0] ramaddrext=6'b000000;			// RAM address extension 4M RAM (Hannes/Csory)
reg romconfig=0;								// ROM config mode enables a special kernal to configure ROM versions
reg romconfreset=0;
reg [7:0] romreg_data=8'hff;
reg [7:0] plus4_datalatch=8'h0;
reg sreset=1'b1;
reg [23:0] resetcounter=24'b0;
reg [15:0] plus4_addrlatch=16'b0;
wire keyreset;
wire key_esc;
wire [4:0] joy0port,joy1port;				// keyboard emulated joystick ports
wire [4:0] joy0emu,joy1emu;				// keyboard emulated joystick ports masked by select lines 
wire RAS;
wire CAS;
wire RW;
wire cs0;
wire cs1;
wire [35:0] CONTROL0;
wire [3:0] cycle;
reg pla_arm;

wire boot_cs0;
wire boot_cs1;
wire boot_rw;
wire boot_done;
wire cfg_done;
wire sdram_cs0;
wire sdram_cs1;
wire sdram_rw;
wire sdram_cas;
wire [15:0] ram_addr;
wire [5:0] sdram_addrext;
wire [7:0] sdram_datain;
wire flash_clken;
wire trigger;


	
// Instantiate the clock module, produce 28.375 Mhz clock for PAL Plus4
palclockgen PAL_PLL
   (// Clock in ports
    .CLK_IN1(CLK32),      					// Papilio Pro platform's clock in
    // Clock out ports
    .CLK_OUT1(CLK28)     					// 28 Mhz clock
    // Status and control signals
    );       // IN


// Generate SDRAM clock signal. It provides a 180 degree shifted clk from FPGA global clock
// The module used here is Xilinx specific, for other FPGA vendors use different method to generate SDRAM_CLK
// See FPGA documentation on how to generate a clock signal on a user IO pin
	sdram_clk ram_clk (
		.clk(CLK28),
		.sdram_clk(SDRAM_CLK)
		);

// 8501 CPU
/*	mos8501 cpu (							// 8501 using FPGA64 cpu core
		.clk(CLK28), 
		.reset(sreset), 
		.enable(cpuenable),  
		.irq_n(irq_n), 
		.data_in(plus4_data), 
		.data_out(cpu_data), 
		.address(cpu_addr),
		.gate_in(mux),
		.rw(RW),								// rw=high read, rw=low write
		.port_in(port_in),
		.port_out(port_out),
		.rdy(rdy),
		.aec(aec)
	); */
	
mos8501_t65 cpu (							// 8501 using T65 core
		.clk(CLK28), 
		.reset(sreset), 
		.enable(cpuenable),  
		.irq_n(irq_n), 
		.data_in(plus4_data), 
		.data_out(cpu_data), 
		.address(cpu_addr),
		.gate_in(mux),
		.rw(RW),								// rw=high read, rw=low write
		.port_in(port_in),
		.port_out(port_out),
		.rdy(rdy),
		.aec(aec)
);

// TED 8360 instance	

ted mos8360(
	.clk(CLK28),
	.addr_in(plus4_addr),
	.addr_out(ted_addr),
	.data_in(plus4_data),
	.data_out(ted_data),
	.rw(RW),
	.cpuclk(phi0),							// phi0 is used for a real external 8501 CPU and internal/external PLA
	.color(plus4_color),
	.csync(HSYNC),
	.irq(irq_n),
	.ba(rdy),
	.mux(mux),
	.ras(RAS),
	.cas(CAS),
	.cs0(cs0),
	.cs1(cs1),
	.aec(aec),
	.k(kbus),
	.snd(sound),
	.cpuenable(cpuenable),
	.pal()
	);

// SDRAM controller
 sdram_controller ram_ctrl(
		.sdram_addr(SDRAM_ADDR),
		.sdram_data(SDRAM_DATA),
		.sdram_dqm({SDRAM_DQMH,SDRAM_DQML}),
		.sdram_ba(SDRAM_BA),
		.sdram_we(SDRAM_nWE),
		.sdram_ras(SDRAM_nRAS),
		.sdram_cas(SDRAM_nCAS),
		.sdram_cs(SDRAM_CS),
		.sdram_cke(SDRAM_CKE),
		.clk(CLK28),
		.plus4_addr(ram_addr),
		.plus4_addrext(sdram_addrext),								
		.plus4_ras(RAS),
		.plus4_cas(sdram_cas),
		.plus4_rw(sdram_rw),
		.plus4_cs0(sdram_cs0),
		.plus4_cs1(sdram_cs1),
		.ram_datain(sdram_datain),
		.ram_dataout(ram_data),
		.initdone(raminitdone)
 );

// SDRAM connection multiplexers

assign ram_addr=(cfg_done)?plus4_addr:boot_addr;
assign sdram_addrext=(boot_done)?plus4_addrext:boot_addrext;
assign sdram_cs0=(boot_done)?cs0:boot_cs0;
assign sdram_cs1=(boot_done)?cs1:boot_cs1;
assign sdram_rw=(boot_done)?RW:boot_rw;
assign sdram_datain=(boot_done)?plus4_data:boot_data;
assign sdram_cas=(boot_done)?CAS:1'b1;

assign plus4_addrext=(~cs0|~cs1)?romaddrext:ramaddrext;	// set ROM or RAM address extension


// Color decoder to 12bit RGB	
 
colors_to_rgb colordecode (
	.clk(CLK28),
	.color(plus4_color),
	.red(RED),
	.green(GREEN),
	.blue(BLUE)
	);

// keyboard part

ps2receiver ps2rcv(
    .clk(CLK28),
    .ps2_clk(PS2CLK),
    .ps2_data(PS2DAT),
    .rx_done(keyreceived),
    .ps2scancode(keyscancode)
    );

c16_keymatrix keyboard(
	 .clk(CLK28),
    .scancode(keyscancode),
    .receiveflag(keyreceived),
	 .row(keyboard_row),
    .kbus(key),
	 .keyreset(keyreset),
	 .joy0(joy0port),
	 .joy1(joy1port),
	 .esc(key_esc)
    );

mos6529 keyport(
	 .clk(CLK28),
    .data_in(plus4_data),
    .data_out(keyport_data),
    .port_in(keyboard_row),	// keyport 6529 in C16/Plus4 is unidirectional however if we read it the last written data is read back so we feed back its output.
    .port_out(keyboard_row),
    .rw(RW),
    .cs(FD3x)
    );

// Bootstrap uploads ROM images and CFG registers from Papilio Pro board's SPI flash chip to SDRAM

 bootstrap boot(
	// SPI flash signals
    .flash_cs(FLASH_CS),
	 .flash_ck(FLASH_CK),
	 .flash_si(FLASH_SI),
	 .flash_so(FLASH_SO),
	// generated ROM signals
	 .cs0(boot_cs0),
	 .cs1(boot_cs1),
	 .rw_out(boot_rw),
	 .addr_out(boot_addr),				
	 .addr_ext(boot_addrext),
	 .data_out(boot_data),
	 
	 .reset(1'b0),
	 .boot_enable(raminitdone),
	 .boot_done(boot_done),
	 .cfg_done(cfg_done),
	 .phi(phi0),
	 .clk(CLK28),
	 // signals for SPI FLASH communication via Plus4 bus
	 .cs(boot_cs),
	 .rw_in(RW),
	 .data_in(plus4_data),
	 .addr_in(plus4_addr[2:0])
    );


	
assign AUDIO_R=sound;
assign AUDIO_L=sound;
assign VSYNC=1'b1;										// set scart mode to RGB for TV

// PLA functions derived from TED System Hardware Manual equation table

always @(posedge CLK28) begin							// arm function needs to be registered
	pla_arm<=mux|(~RAS&phi0&pla_arm);
	end

assign KERN=(plus4_addr[15:8]==8'hfc)?1'b1:1'b0;
assign FD3x=((plus4_addr[15:4]==12'hfd3) & pla_arm & phi0 & ~RAS)?1'b1:1'b0;	// KEYPORT
assign FDDx=((plus4_addr[15:4]==12'hfdd) & pla_arm & phi0 & ~RAS)?1'b1:1'b0;	// ADDR CLK
assign FD0x=((plus4_addr[15:4]==12'hfd0) & phi0)?1'b1:1'b0;  						// 6551
assign FD1x=((plus4_addr[15:4]==12'hfd1) & pla_arm & phi0 & ~RAS)?1'b1:1'b0;  // 6529
assign phi2=~RAS & pla_arm & phi0;															// PHI2 CLK not used at the moment
assign FD2x=((plus4_addr[15:4]==12'hfd2) & phi0 & ~RAS); 							//SPEECH $FD2X is not used in Plus4 (used for Commodore 364)
assign FD9x=((plus4_addr[15:4]==12'hfd9) & phi0 & ~RAS);								// FPGATED configuration register

// ROM MMU 

always @(posedge CLK28) begin									// Plus4 motherboard ROM selector register (U21)
	FDDx_prev<=FDDx;
	if(sreset)
		romselect<=4'h0;
	else if(~FDDx_prev & FDDx & ~RW)
		romselect<=plus4_addr[3:0];
end

always @*	begin													// generating ROM address extension for different ROM versions
		if(~cs0) begin												// low ROM
			case(romselect[1:0])									// based on romselect register set romversion to the active rom version (version 1-16)
					2'b00:	romversion=Basicver;				
					2'b01:	romversion=FunctionLver;
					2'b10:	romversion=C1Lver;
					2'b11:	romversion=C2Lver;
			endcase
			romaddrext={romversion,romselect[1:0]};
		end
		else begin													// high ROM
				case(romselect[3:2])
					2'b00:	romversion=Kernalver;
					2'b01:	romversion=FunctionHver;
					2'b10:	romversion=C1Hver;
					2'b11:	romversion=C2Hver;
				endcase	
				romaddrext=(romconfig)?{4'hf,2'b00}:(KERN)?{Kernalver,2'b00}:{romversion,romselect[3:2]};
		end
end

// ROM config mode flag

always @(posedge CLK28)
	begin
	if(sreset&key_esc)					// activate ROM configuration mode when ESC key is pressed during bootstrap
		romconfig<=1'b1;
	else if(sreset)						// inactivate ROM configuration mode at beginning of hard reset
		romconfig<=1'b0;
	end

// FPGATED ROM config register  (could be placed to a separate module)

always @(posedge CLK28)
	begin
	FD9x_prev<=FD9x;
	phi0_prev<=phi0;
	end


always @(posedge CLK28) begin
	romreg_data<=8'hff;
	romconfreset<=1'b0;
	if(FD9x & RW) begin																// ROM and FPGATED config registers read					
			case(plus4_addr[3:0])
				4'h0:	romreg_data<={Kernalver,Basicver};
				4'h1:	romreg_data<={FunctionHver,FunctionLver};
				4'h2:	romreg_data<={C1Hver,C1Lver};
				4'h3:	romreg_data<={C2Hver,C2Lver};
				default:romreg_data<=8'hff;
			endcase
		end
	// ROM and FPGATED config registers write (only allowed when RomConfig mode is enabled)
	// this part is connected to bootstrap data and address buses during FPGATED configuration in order to load initial values
	// during normal operation it is connected to Plus4 data and address buses so it can be modified via Plus4 bus cycles
	else if((FD9x_prev & ~FD9x & ~RW & romconfig) || (boot_done & ~cfg_done & phi0_prev & ~phi0 & ~boot_rw ))
		begin		
			case(ram_addr[3:0])														// ram_addr is boot_addr during bootstrap, plus4_address after FPGTAED is configured
				4'h0: begin
						Kernalver<=config_data[7:4];								// config_data is boot_data during bootstrap, plus4_datalatch after FPGATED is configured
						Basicver<=config_data[3:0];
						end
				4'h1:	begin
						FunctionHver<=config_data[7:4];
						FunctionLver<=config_data[3:0];
						end
				4'h2:	begin
						C1Hver<=config_data[7:4];
						C1Lver<=config_data[3:0];
						end
				4'h3:	begin
						C2Hver<=config_data[7:4];
						C2Lver<=config_data[3:0];
						end
				4'h4: begin														// Config register 1
				// add config register write here
						end
				4'h5:	begin														// Config register 2
				// add config register write here
						end
				4'h7: begin
						romconfreset<=1'b1;									// Reset system when writing to this address
						end
			endcase
		end
end

assign boot_cs=FD9x&plus4_addr[3]&(~cfg_done|romconfig);			// FPGATED boot chipselect signal 
assign config_data=(cfg_done)?plus4_datalatch:boot_data; 			// data for config registers write is taken from Plus4 databus or boot databus

// Plus4 reset circuit

always @(posedge CLK28)		// reset tries to emulate the length of a real reset
	begin
	if(RESET|keyreset|romconfreset)		// reset can be triggered by reset button , CTRL+ALT+DEL from keyboard or from ROM config kernal
		begin
		resetcounter<=0;		// start reset length counter
		sreset<=1;				// set synchronous reset for CPU
		end
	else begin
		if(resetcounter==24'd16777215) begin
			if(boot_done & cfg_done)
				sreset<=0;			// end of reset after approximately 590ms
			end
		else begin
			resetcounter<=resetcounter+24'b1;
			sreset<=1;
			end
		end
	end	

	
// Motherboard bus connections

assign plus4_addr=(~mux)?plus4_addrlatch:cpu_addr&ted_addr;																					// Plus4 address bus
assign plus4_data=(mux)?plus4_datalatch:cpu_data&ted_data&ram_data&keyport_data&romreg_data&boot_data;						// Plus4 data bus using sdram for ROM

always @(posedge CLK28)							// address and data bus latching emulates dynamic memory behaviour of these buses 
	begin
	plus4_datalatch<=plus4_data;
	plus4_addrlatch<=plus4_addr;
	end

// Joystick and Keyboard connection to keybus

assign joy0emu=(~plus4_data[2])?joy0port:5'b11111;			// keyboard emulated joy0 port is allowed to kbus only when its select line is active (D2 bit)
assign joy1emu=(~plus4_data[1])?joy1port:5'b11111;			// keyboard emulated joy1 port is allowed to kbus only when its select line is active (D1 bit)

assign kbus={key[7]&joy1emu[4],key[6]&joy0emu[4],key[5:4],key[3]&joy0emu[3]&joy1emu[3],key[2]&joy0emu[2]&joy1emu[2],key[1]&joy0emu[1]&joy1emu[1],key[0]&joy0emu[0]&joy1emu[0]};

// connect IEC bus

assign IEC_DATAOUT=port_out[0];
assign port_in[7]=IEC_DATAIN;
assign IEC_CLKOUT=port_out[1];
assign port_in[6]=IEC_CLKIN;
assign IEC_ATNOUT=port_out[2];
//assign ATN=IEC_ATNIN;
assign IEC_RESET=sreset;


chipscope_icon plus4_ICON (
    .CONTROL0(CONTROL0) // INOUT BUS [35:0]
);
chipscope_ila plus4_ILA (
    .CONTROL(CONTROL0), // INOUT BUS [35:0]
    .CLK(CLK28), // IN
//    .TRIG0({trigger,FLASH_CS,flash_clken,FLASH_SI,FLASH_SO,boot_cs0,boot_cs1,boot_rw,boot_addr,boot_addrext,boot_data,phi0,begin_boot}) // IN BUS [39:0]
	.TRIG0({plus4_addr,plus4_data}), // IN BUS [23:0]
	.TRIG1({sreset,romconfig,irq_n,phi0,RW,romaddrext,cs0,cs1,mux,aec,rdy}) // IN BUS [15:0]
);

endmodule
